----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    01:54:34 06/02/2011 
-- Design Name: 
-- Module Name:    sha256_s0 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity sha256_s0 is
    Port ( d : in  STD_LOGIC_VECTOR (31 downto 0);
           q : out  STD_LOGIC_VECTOR (31 downto 0));
end sha256_s0;

architecture Behavioral of sha256_s0 is

begin

	q(31 downto 29) <= d(6 downto 4) xor d(17 downto 15);
	q(28 downto 0) <= (d(3 downto 0) & d(31 downto 7)) xor (d(14 downto 0) & d(31 downto 18)) xor d(31 downto 3);

end Behavioral;

